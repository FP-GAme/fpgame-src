module vram_rd_sel (

);

endmodule : vram_rd_sel
