module vram_sync_writer (

    // from vram 1
    output logic [] pram1_addr,
    input  logic [] pram1_rddata,
    input  logic [] pram2_wrdata,

    // from vram 2

);



endmodule : vram_sync_writer
