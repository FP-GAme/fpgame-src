module row_ram_swap (
    input  logic clk,
    input  logic rst_n,

    // From/to hdmi_video_output (reader)
    input  logic        rowram_swap,
    output logic [9:0]  hdmi_rowram_rddata,
    input  logic [8:0]  hdmi_rowram_rdaddr,

    // From Pixel Mixer (writer)
    input  logic [9:0]  pmxr_rowram_wrdata,
    input  logic [8:0]  pmxr_rowram_wraddr,
    input  logic        pmxr_rowram_wren
);
    // Flip-Flop to store swapped state after the rowram_swap signal is received.
    logic swapped;

    // Every time we see the swap signal, we need to ignore the next time we see it.
    // This is because the swap signal is generated by a 25MHz clock, and we are running a 50MHz
    //   clock: Our 50MHz clock effectively sees 2 25MHz clocks worth of that swap signal.
    logic ignore_swap;

    logic [8:0] rr1_addr,   rr2_addr;
    logic [9:0] rr1_rddata, rr2_rddata;
    logic [9:0] rr1_wrdata, rr2_wrdata;
    logic       rr1_wren,   rr2_wren;

    // TODO REMOVE AFTER DEBUG:
    // THIS WORKED
    /*row_ram rr1 (
        .address_a(hdmi_rowram_rdaddr),
        .address_b(9'b0),
        .clock(clk),
        .data_a(10'b0), // TODO Change
        .data_b(10'b0), // TODO Change
        .wren_a(1'b0), // TODO Change
        .wren_b(1'b0), // TODO Change
        .q_a(hdmi_rowram_rddata),
        .q_b()
    );*/

    // Even though we have dual-ports, we simplify things by using 1 port (ignoring port b)
    row_ram rr1 (
        .address_a(rr1_addr),
        .address_b(9'b0),
        .clock(clk),
        .data_a(rr1_wrdata),
        .data_b(10'b0),
        .wren_a(rr1_wren),
        .wren_b(1'b0),
        .q_a(rr1_rddata),
        .q_b()
    );
    row_ram rr2 (
        .address_a(rr2_addr),
        .address_b(9'b0),
        .clock(clk),
        .data_a(rr2_wrdata),
        .data_b(10'b0),
        .wren_a(rr2_wren),
        .wren_b(1'b0),
        .q_a(rr2_rddata),
        .q_b()
    );

    // The default state (rowram_swapped=0):
    //   hdmi_video_output rd rr1
    //   pixel_mixer       wr rr2
    // The swapped state (rowram_swapped=1):
    //   hdmi_video_output rd rr2
    //   pixel_mixer       wr rr1

    assign rr1_addr = (swapped) ? pmxr_rowram_wraddr : hdmi_rowram_rdaddr;
    assign rr1_wren = (swapped) ? pmxr_rowram_wren : 1'b0;
    // wrdata is safe to tie to both RAMs. It is essentially a "don't-care", so the wren must be 0
    //   on the RAM we don't intend on writing to. This RAM not being written to is, of course,
    //   being read by the hdmi_video_output, so this should be safe by default.
    // TODO: Unlikely, but if necessary, use actual don't-cares. Increases complexity but may improve timing.
    assign rr1_wrdata = pmxr_rowram_wrdata;

    assign rr2_addr = (swapped) ? hdmi_rowram_rdaddr : pmxr_rowram_wraddr;
    assign rr2_wren = (swapped) ? 1'b0 : pmxr_rowram_wren;
    assign rr2_wrdata = pmxr_rowram_wrdata;

    assign hdmi_rowram_rddata = (swapped) ? rr2_rddata : rr1_rddata;

    /*assign rr1_addr = hdmi_rowram_rdaddr;
    assign hdmi_rowram_rddata = rr1_rddata;
    assign rr1_wren = 1'b0;
    assign rr1_wrdata = 10'b0;*/

    // Receive buffer swap signal. Buffers are swapped combinationally after the clock edge after
    //   the rowram_swap signal has been detected.
    always_ff @(posedge clk, negedge rst_n) begin
        if (!rst_n) begin
            swapped <= 1'b0;
            ignore_swap <= 1'b0;
        end
        else if (rowram_swap) begin
            //swapped <= 1'b0; // TODO: Remove after debug
            //ignore_swap <= 1'b0; // TODO: Remove after debug
            swapped <= (ignore_swap) ? swapped : ~swapped;
            ignore_swap <= ~ignore_swap;
        end
    end
endmodule : row_ram_swap