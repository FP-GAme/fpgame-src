module ppu (

);

endmodule : ppu
